library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity cajitaAnds is
port
(
	entradaZeroAlu, entradaBranch, entradaPcWrite : in std_logic;
	senalSalida : out std_logic
);

end cajitaAnds;

architecture arch of cajitaAnds is
begin
	process (entradaZeroAlu, entradaBranch, entradaPcWrite)
	begin
		senalSalida <= (entradaZeroAlu and entradaBranch) or entradaPcWrite;
	end process;
end arch;